`timescale 1ns / 1ps
`include "config.v"

module mem_ctrl